`include "wr_xtn.sv"
`include "my_sequence.sv"
`include "my_reset_sequence.sv"
`include "my_driver_callback.sv"

`include "my_wr_sequencer.sv"
`include "my_wr_driver.sv"
`include "my_wr_monitor.sv"

`include "my_wr_agent.sv"
`include "my_env.sv"
`include "base_test.sv"